module bloodAbnormalityDetector(
 bloodPH,
 bloodType,
 bloodAbnormality);
input [3:0] bloodPH;
input [2:0] bloodType;
output bloodAbnormality;
 // write your code here, please.
endmodule
