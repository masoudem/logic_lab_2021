module temperatureAbnormalityDetector(
 bloodSensor,
 glycemicIndex);
input [7:0] bloodSensor;
output [3:0] glycemicIndex;
 // write your code here, please.
endmodule
