/*--  *******************************************************
--  Computer Architecture Course, Laboratory Sources 
--  Amirkabir University of Technology (Tehran Polytechnic)
--  Department of Computer Engineering (CE-AUT)
--  https://ce[dot]aut[dot]ac[dot]ir
--  *******************************************************
--  All Rights reserved (C) 2020-2021
--  *******************************************************
--  Student ID  : 
--  Student Name: 
--  Student Mail: 
--  *******************************************************
--  Additional Comments:
--
--*/

/*-----------------------------------------------------------
---  Module Name: bfpfemale
-----------------------------------------------------------*/
`timescale 1 ns/1 ns
module bfpfemale(
w,
h,
a,
bfprange);
  input [7:0] w;
  input [7:0] h;
  input [7:0] a;
  output [7:0] range;
 // write your code here, please.
endmodule
