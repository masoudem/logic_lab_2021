module temperatureAbnormalityDetector(
 factotyBaseTemp,
 factotyTempCoef,
 tempSensorValue,
 temperatureAbnormality);
input [4:0] factotyBaseTemp;
input [3:0] factotyTempCoef;
input [3:0] tempSensorValue;
output temperatureAbnormality;
 // write your code here, please.
endmodule
