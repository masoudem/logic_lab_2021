module pressureAbnormalityDetector(
 pressureData,
 presureAbnormality);
input [5:0] pressureData;
output presureAbnormality;
 // write your code here, please.
endmodule
