module fallingDetector(
 fdSensorValue,
 fdFactoryValue,
 fallDetected);
input [7:0] fdSensorValue;
input [7:0] fdFactoryValue;
output fallDetected;
 // write your code here, please.
endmodul
