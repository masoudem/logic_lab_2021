/*--  *******************************************************
--  Computer Architecture Course, Laboratory Sources 
--  Amirkabir University of Technology (Tehran Polytechnic)
--  Department of Computer Engineering (CE-AUT)
--  https://ce[dot]aut[dot]ac[dot]ir
--  *******************************************************
--  All Rights reserved (C) 2020-2021
--  *******************************************************
--  Student ID  : 
--  Student Name: 
--  Student Mail: 
--  *******************************************************
--  Additional Comments:
--
--*/

/*-----------------------------------------------------------
---  Module Name: bloodPHAnalyzer
-----------------------------------------------------------*/
`timescale 1 ns/1 ns
module bloodPHAnalyzer(
 bloodPH,
 abnormalityP,
 abnormalityQ);
input [3:0] bloodPH;
output abnormalityP;
output abnormalityQ;
 // write your code here, please.
endmodule
