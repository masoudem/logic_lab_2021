module pressureAnalyzer(
 pData,
 pWarning);
input [4:0] pData;
output pDarning;
 // write your code here, please.
endmodule
