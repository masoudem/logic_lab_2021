module bloodPHAnalyzer(
 bloodPH,
 abnormalityP,
 abnormalityQ);
input [3:0] bloodPH;
output abnormalityP;
output abnormalityQ;
 // write your code here, please.
endmodule
