/*--  *******************************************************
--  Computer Architecture Course, Laboratory Sources 
--  Amirkabir University of Technology (Tehran Polytechnic)
--  Department of Computer Engineering (CE-AUT)
--  https://ce[dot]aut[dot]ac[dot]ir
--  *******************************************************
--  All Rights reserved (C) 2020-2021
--  *******************************************************
--  Student ID  : 
--  Student Name: 
--  Student Mail: 
--  *******************************************************
--  Additional Comments:
--
--*/

/*-----------------------------------------------------------
---  Module Name: bfpmale
-----------------------------------------------------------*/
`timescale 1 ns/1 ns
module bfpmale(
wm,
hm,
am,
bfprange);
  input [7:0] wm;
  input [7:0] hm;
  input [7:0] am;
  output [7:0] rangem;
 // write your code here, please.
endmodule
