/*--  *******************************************************
--  Computer Architecture Course, Laboratory Sources 
--  Amirkabir University of Technology (Tehran Polytechnic)
--  Department of Computer Engineering (CE-AUT)
--  https://ce[dot]aut[dot]ac[dot]ir
--  *******************************************************
--  All Rights reserved (C) 2020-2021
--  *******************************************************
--  Student ID  : 
--  Student Name: 
--  Student Mail: 
--  *******************************************************
--  Additional Comments:
--
--*/

/*-----------------------------------------------------------
---  Module Name: bmd 
-----------------------------------------------------------*/
`timescale 1 ns/1 ns
module bfpfemale(
bmdrange,
normal,
abnormal);
  input [1:0] bmdrange;
  output normal;
  output abnormal;
 // write your code here, please.
endmodule
