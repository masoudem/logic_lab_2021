module parityErrorChecker(
 data,
 error);
input [5:0] data;
output error;
 // write your code here, please.
endmodule
