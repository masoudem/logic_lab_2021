module temperatureCalculator(
 factotyBaseTemp,
 factotyTempCoef,
 tempSensorValue,
 temperature);
input [4:0] factotyBaseTemp;
input [3:0] factotyTempCoef;
input [3:0] tempSensorValue;
output [7:0] temperature;
 // write your code here, please.
endmodule
