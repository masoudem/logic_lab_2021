/*--  *******************************************************
--  Computer Architecture Course, Laboratory Sources 
--  Amirkabir University of Technology (Tehran Polytechnic)
--  Department of Computer Engineering (CE-AUT)
--  https://ce[dot]aut[dot]ac[dot]ir
--  *******************************************************
--  All Rights reserved (C) 2020-2021
--  *******************************************************
--  Student ID  : 
--  Student Name: 
--  Student Mail: 
--  *******************************************************
--  Additional Comments:
--
--*/

/*-----------------------------------------------------------
---  Module Name: bloodTypeClassification 
-----------------------------------------------------------*/
`timescale 1 ns/1 ns
module bloodTypeClassification(
 bloodType,
 bloodClass);
input [2:0] bloodType;
output bloodClass;
 // write your code here, please.
endmodule
