/*--  *******************************************************
--  Computer Architecture Course, Laboratory Sources 
--  Amirkabir University of Technology (Tehran Polytechnic)
--  Department of Computer Engineering (CE-AUT)
--  https://ce[dot]aut[dot]ac[dot]ir
--  *******************************************************
--  All Rights reserved (C) 2020-2021
--  *******************************************************
--  Student ID  : 
--  Student Name: 
--  Student Mail: 
--  *******************************************************
--  Additional Comments:
--
--*/

/*-----------------------------------------------------------
---  Module Name: bfpfemale
-----------------------------------------------------------*/
`timescale 1 ns/1 ns
module bfpfemale(
w,
h,
a,
bfprange);
  input [7:0] wf;
  input [7:0] hf;
  input [7:0] af;
  output [7:0] rangef;
 // write your code here, please.
endmodule
