`timescale 1ns / 1ps
/*--  *******************************************************
--  Computer Architecture Course, Laboratory Sources 
--  Amirkabir University of Technology (Tehran Polytechnic)
--  Department of Computer Engineering (CE-AUT)
--  https://ce[dot]aut[dot]ac[dot]ir
--  *******************************************************
--  All Rights reserved (C) 2021-2022
--  *******************************************************
--  Student ID  : 
--  Student Name: 
--  Student Mail: 
--  *******************************************************
--  Additional Comments:
--
--*/

/*-----------------------------------------------------------
---  Module Name: controller_and_register
-----------------------------------------------------------*/

module controller_and_register(confirm, request, clock, inputData, dataQ, dataP);
input confirm, request, clock;
input [7:0] inputData;
output [6:0] dataQ, dataP;
 // write your code here, please.
endmodule
